///////////////////////////////////////////////////////////////////////////////
// File       : riscv_top.sv
// Ver        : 0.1
// Date       : 06.01.2024
///////////////////////////////////////////////////////////////////////////////
//
// Description: This is my 5-stage pipeline implementation of cv32e40p equivalent
//
///////////////////////////////////////////////////////////////////////////////
//
// Authors    : Yunhai Qiao (dellysunny@yahoo.com)
//
///////////////////////////////////////////////////////////////////////////////

